library verilog;
use verilog.vl_types.all;
entity bcd_7seg_vlg_vec_tst is
end bcd_7seg_vlg_vec_tst;
